`timescale 1 ns / 1 ps

module adc_test_streamer_v2_0_M00_AXIS #
(
    // Users to add parameters here

    // User parameters ends

    parameter integer C_M_AXIS_TDATA_WIDTH	= 64,
    // Start count is the number of clock cycles the master will wait before initiating/issuing any transaction.
    parameter integer C_M_START_COUNT	= 32
)
(
    // Users to add ports here
    input wire [63:0] ADC_BUS,
    input wire ADC_DATA_CLK,
    input wire ADC_DATA_VALID,
    input wire ADC_FIFO_RESET,
    input wire ADC_EOF,
    
    output wire [5:0] dbg_adcstream_state,
    output wire dbg_axi_rdy,
    output wire dbg_acq_axi_running,
    output wire [31:0] dbg_acq_axi_upcounter,
    output wire [31:0] dbg_acq_axi_downcounter,
    output wire [10:0] dbg_acq_trigger_out_ctr,
    output wire [15:0] dbg_rd_data_count,
    output wire [15:0] dbg_wr_data_count,

    input ACQ_RUN,
    input ACQ_ABORT,
    input ACQ_TRIG_MASK,
    input ACQ_TRIG_RST,
    input ACQ_DEPTH_MUX,
    input [28:0] ACQ_DEPTH_A,
    input [28:0] ACQ_DEPTH_B,
    output reg ACQ_DONE,
    output reg ACQ_HAVE_TRIG,
    input ACQ_AXI_RUN,
    output ACQ_FULL_DATA_LOSS,
    
    input TRIGGER_IN,
    output reg TRIGGER_OUT,
    output reg [31:0] TRIGGER_POS,
    input [2:0] TRIGGER_SUB_WORD,
    
    // User ports ends
    // Do not modify the ports beyond this line

    // Global ports
    input wire  M_AXIS_ACLK,
    // 
    input wire  M_AXIS_ARESETN,
    // Master Stream Ports. TVALID indicates that the master is driving a valid transfer, A transfer takes place when both TVALID and TREADY are asserted. 
    output wire  M_AXIS_TVALID,
    // TDATA is the primary payload that is used to provide the data that is passing across the interface from the master.
    output wire [C_M_AXIS_TDATA_WIDTH-1 : 0] M_AXIS_TDATA,
    // TSTRB is the byte qualifier that indicates whether the content of the associated byte of TDATA is processed as a data byte or a position byte.
    output wire [(C_M_AXIS_TDATA_WIDTH/8)-1 : 0] M_AXIS_TSTRB,
    // TLAST indicates the boundary of a packet.
    output wire  M_AXIS_TLAST,
    // TREADY indicates that the slave can accept a transfer in the current cycle.
    input wire  M_AXIS_TREADY
);               
                                                                           
parameter ST_IDLE = 0;                                                               
parameter ST_STREAMING = 1;                                                          
parameter ST_STOP_TRIGGERED = 2;                                                     
parameter ST_STOP_EOF = 3;

// Debug signals
assign dbg_axi_rdy = M_AXIS_TREADY;
assign dbg_acq_axi_running = acq_axi_running;
assign dbg_adcstream_state = adcstream_state;
assign dbg_trigger_out_ctr = trigger_out_ctr;
assign dbg_acq_axi_upcounter = acq_axi_upcounter;
assign dbg_acq_axi_downcounter = acq_axi_downcounter;
assign dbg_acq_trigger_out_ctr = dbg_acq_trigger_out_ctr;

reg [5:0] adcstream_state = ST_IDLE;

reg acq_tvalid = 0;
reg acq_axi_running = 0;

reg acq_gen_tlast = 0; 
reg acq_gen_tvalid_mask = 0;
reg [1:0] acq_gen_tlast_ctr = 0;
 
reg [10:0] trigger_out_ctr;

// TODO: try to figure out how we could common these counters
reg [28:0] acq_axi_downcounter = 0;
reg [28:0] acq_axi_upcounter = 0;

wire [63:0] fifo_data_out;

reg adc_fifo_full_latch = 0;
assign ACQ_FULL_DATA_LOSS = adc_fifo_full_latch;

// TVALID is high when: FIFO reset not busy,  FIFO not almost empty
assign M_AXIS_TVALID = /*(!fifo_rd_busy) && */(!fifo_almost_empty) && acq_gen_tvalid_mask; 
assign M_AXIS_TDATA	= fifo_data_out;
assign M_AXIS_TLAST	= acq_gen_tlast; 

// TSTRB == not used (set to all 1's)
assign M_AXIS_TSTRB	= {(C_M_AXIS_TDATA_WIDTH/8){1'b1}};

wire fifo_almost_empty;
wire fifo_full;

// Output busy signals from the FIFO generator
wire fifo_wr_busy;
wire fifo_rd_busy;

// Write enabled when ADC_VALID asserted (Data should start filling FIFO; DMA will ready when ready)
wire fifo_wr_en = ADC_DATA_VALID;                             
 
// Read enabled when TREADY asserted & data available in FIFO & acq_axi_running asserted & TVALID present
wire fifo_rd_en = M_AXIS_TREADY && (!fifo_almost_empty) && acq_axi_running && acq_gen_tvalid_mask;        

// FIFO reset a combination of AXI reset and external slow reset signal
wire fifo_int_reset = ((!M_AXIS_ARESETN) || ADC_FIFO_RESET);    

// FIFO data in and data out consists of trigger_signal + 64-bit data.  
wire [64:0] fifo_data_in = {(TRIGGER_IN && !ACQ_TRIG_MASK), ADC_BUS};
wire [64:0] fifo_data_out;

assign fifo_out_trigger = fifo_data_out[64];

// FIFO generator connection (block design)
fifo_generator_0 fifo_generator_0_inst (
    .full(ADC_FIFO_FULL),
    .wr_en(fifo_wr_en),
    .prog_empty(fifo_almost_empty),
    .rd_en(fifo_rd_en),
    .din(fifo_data_in),
    .wr_clk(ADC_DATA_CLK),
    .dout(fifo_data_out),
    .rd_clk(M_AXIS_ACLK),
    .rst(fifo_int_reset),
    .rd_data_count(dbg_rd_data_count),
    .wr_data_count(dbg_wr_data_count)
    //.wr_rst_busy(fifo_wr_busy),
    //.rd_rst_busy(fifo_rd_busy)
);

/*
 * State machine.  This runs on the AXI bus clock. 
 */
always @(posedge M_AXIS_ACLK) begin

    /*
     * Trigger out generator.  Generate a 16-clock pulse every time a trigger
     * is accepted by the acquisition engine.  Note this is NOT the same as 
     * the direct trigger signal.  Also note the output pulse width is a multiple
     * of the AXI bus clock, which should be fixed by design.
     */
    if (trigger_out_ctr > 1) begin
        trigger_out_ctr <= trigger_out_ctr - 1;
        TRIGGER_OUT <= 1;
    end else begin
        TRIGGER_OUT <= 0;
    end
    
    /*
     * If FIFO_FULL goes high then we set a state which is only cleared by starting
     * a new acquisition.  This signal indicates data has been lost and the FIFO must
     * be reset to avoid data corruption.
     */
    if (ADC_FIFO_FULL) begin
        adc_fifo_full_latch <= 1;
    end

    case (adcstream_state) 
    
        ST_IDLE : begin
            if (ACQ_AXI_RUN && M_AXIS_TREADY) begin
                ACQ_HAVE_TRIG <= 0;
                ACQ_DONE <= 0;
                
                // Load the required downcounter
                if (!ACQ_DEPTH_MUX) begin
                    acq_axi_downcounter <= ACQ_DEPTH_A;
                end else begin
                    acq_axi_downcounter <= ACQ_DEPTH_B;
                end
                
                acq_axi_upcounter <= 0;
                
                // Invalid TRIGGER_POS:  Acq not yet run
                TRIGGER_POS <= 32'hfffffffe;
                
                adc_fifo_full_latch <= 0;
                acq_axi_running <= 1;
                //adcclkdm_tvalid_init <= 1;
                adcstream_state <= ST_STREAMING;
            end
        end
        
        ST_STREAMING : begin
            // Only adjust counters and handle triggers, etc. if data is available in FIFO.
            if ((!fifo_almost_empty) && M_AXIS_TREADY && (!M_AXIS_TLAST)) begin
                acq_axi_upcounter <= acq_axi_upcounter + 1;
                acq_axi_downcounter <= acq_axi_downcounter - 1;
            
                if (acq_axi_downcounter == 0) begin
                    // Trigger not valid in this instance; set TRIGGER_POS to invalid value
                    adcstream_state <= ST_STOP_EOF;
                    TRIGGER_POS <= 32'hffffffff;
                    
                    // Start TLAST pulse generation. TVALID stays active until 1 cycle of TLAST.
                    acq_gen_tvalid_mask <= 1;
                    acq_gen_tlast <= 1;
                end else if (fifo_out_trigger) begin
                    adcstream_state <= ST_STOP_TRIGGERED;
                    
                    // Start TLAST pulse generation. TVALID stays active until 1 cycle of TLAST.
                    acq_gen_tvalid_mask <= 1;
                    acq_gen_tlast <= 1;
                
                    // Load merged trigger position register (32 bits)
                    TRIGGER_POS <= {2'b00, acq_axi_upcounter, TRIGGER_SUB_WORD};
                    
                    // Load trigger counter to generate trigger pulse (1us at ~177MHz)
                    // TODO: this might be application configurable to consistently generate the same pulse
                    // width at different sample rates, also for user configurability if desired.
                    trigger_out_ctr <= 177; 
                end else begin
                    // Otherwise, assert TVALID while streaming data.
                    acq_gen_tvalid_mask <= 1;
                    acq_gen_tlast <= 0;
                end
            end
        end
        
        ST_STOP_TRIGGERED : begin
            // Leave IOs in the "stopped-with-trig" state;  to exit this state the 
            // PS must drive ACQ_AXI_RUN low
            ACQ_HAVE_TRIG <= 1;
            ACQ_DONE <= 1;
            
            // Stop sending TLAST signal, stop sending VALID signal
            acq_gen_tlast <= 0;
            acq_gen_tvalid_mask <= 0;
                    
            if (!ACQ_AXI_RUN) begin
                adcstream_state <= ST_IDLE;
            end
        end
        
        ST_STOP_EOF : begin
            // Leave IOs in the "stopped-with-no-trig" state;  to exit this state the 
            // PS must drive ACQ_AXI_RUN low
            ACQ_HAVE_TRIG <= 0;
            ACQ_DONE <= 1;
            
            // Stop sending TLAST signal, stop sending VALID signal
            acq_gen_tlast <= 0;
            acq_gen_tvalid_mask <= 0;
            
            if (!ACQ_AXI_RUN) begin
                adcstream_state <= ST_IDLE;
            end
        end
    
    endcase

end

endmodule
